module Key2pxl
	(
		input wire [7:0] key,
		input wire [4:0] i_X, 
		input wire [4:0] i_Y,
		output reg o_one_pixel
	);



localparam n1 = 256'b0000_0000_0000_0000_0000_0011_1100_0000_0000_0011_1100_0000_0000_1111_1100_0000_0000_1111_1100_0000_0000_0011_1100_0000_0000_0011_1100_0000_0000_0011_1100_0000_0000_0011_1100_0000_0000_0011_1100_0000_0000_0011_1100_0000_0000_0011_1100_0000_0000_0011_1100_0000_0000_1111_1111_0000_0000_1111_1111_0000_0000_0000_0000_0000;

localparam n2 = 256'b0000_0000_0000_0000_0000_1111_1111_0000_0011_1111_1111_1000_0111_1100_0011_1100_0110_0000_0011_1100_0000_0000_0011_1100_0000_0000_0011_1100_0000_0011_1111_0000_0000_0011_1111_0000_0000_1111_0000_0000_0000_1111_0000_0000_0011_1100_0000_0000_0011_1100_0000_0000_0111_1111_1111_1110_0111_1111_1111_1110_0000_0000_0000_0000;

localparam n3 = 256'b0000_0000_0000_0000_0001_1111_1111_1000_0011_1111_1111_1000_0000_0000_0011_1100_0000_0000_0011_1100_0000_0000_0011_1000_0000_0000_0011_1000_0000_1111_1111_0000_0000_1111_1111_0000_0000_0000_0011_1000_0000_0000_0011_1000_0000_0000_0011_1100_0000_0000_0011_1100_0011_1111_1111_1000_0001_1111_1111_1000_0000_0000_0000_0000;

localparam n4 = 256'b0000_0000_0000_0000_0011_1100_0011_1100_0011_1100_0011_1100_0011_1100_0011_1100_0011_1100_0011_1100_0011_1100_0011_1100_0011_1100_0011_1100_0011_1100_0011_1100_0011_1100_0011_1100_0000_1111_1111_1100_0000_1111_1111_1100_0000_0000_0011_1100_0000_0000_0011_1100_0000_0000_0011_1100_0000_0000_0011_1100_0000_0000_0000_0000;

localparam n5 = 256'b0000_0000_0000_0000_0011_1111_1111_1100_0011_1111_1111_1100_0011_1100_0000_0000_0011_1100_0000_0000_0011_1111_1111_0000_0011_1111_1111_0000_0000_0000_0011_1100_0000_0000_0011_1100_0000_0000_0011_1100_0000_0000_0011_1100_0011_1100_0011_1100_0011_1100_0011_1100_0000_1111_1111_0000_0000_1111_1111_0000_0000_0000_0000_0000;

localparam n6 = 256'b0000_0000_0000_0000_0000_1111_1111_0000_0001_1111_1111_1000_0011_1100_0011_1100_0011_1100_0011_1100_0011_1100_0000_0000_0011_1100_0000_0000_0011_1111_1111_0000_0011_1111_1111_1000_0011_1100_0011_1100_0011_1100_0011_1100_0011_1100_0011_1100_0011_1100_0011_1100_0001_1111_1111_1000_0000_1111_1111_0000_0000_0000_0000_0000;

localparam n7 = 256'b0000_0000_0000_0000_0011_1111_1111_1100_0011_1111_1111_1100_0000_0000_0011_1100_0000_0000_0011_1100_0000_0000_1111_0000_0000_0000_1111_0000_0000_0011_1100_0000_0000_0011_1100_0000_0000_0011_1100_0000_0000_0011_1100_0000_0000_0011_1100_0000_0000_0011_1100_0000_0000_0011_1100_0000_0000_0011_1100_0000_0000_0000_0000_0000;

localparam n8 = 256'b0000_0000_0000_0000_0000_1111_1111_0000_0000_1111_1111_0000_0001_1100_0011_1000_0011_1100_0011_1100_0011_1100_0011_1100_0001_1100_0011_1000_0000_1111_1111_0000_0000_1111_1111_0000_0001_1100_0011_1000_0011_1100_0011_1100_0011_1100_0011_1100_0001_1100_0011_1000_0000_1111_1111_0000_0000_1111_1111_0000_0000_0000_0000_0000;

localparam n9 = 256'b0000_0000_0000_0000_0000_1111_1111_0000_0001_1111_1111_0000_0011_1100_0011_1000_0011_1100_0011_1100_0011_1100_0011_1100_0011_1100_0011_1100_0001_1111_1111_1100_0000_1111_1111_1100_0000_0000_0011_1100_0000_0000_0011_1100_0011_1100_0011_1100_0011_1100_0011_1000_0001_1111_1111_0000_0000_1111_1111_0000_0000_0000_0000_0000;

localparam n0 = 256'b0000_0000_0000_0000_0000_1111_1111_0000_0001_1111_1111_1000_0011_1100_0011_1100_0011_1100_0011_1100_0011_1100_0011_1100_0011_1100_0011_1100_0011_1100_0011_1100_0011_1100_0011_1100_0011_1100_0011_1100_0011_1100_0011_1100_0011_1100_0011_1100_0011_1100_0011_1100_0001_1111_1111_1000_0000_1111_1111_0000_0000_0000_0000_0000;

localparam H =  256'b0000_0000_0000_0000_0011_1000_0001_1100_0011_1000_0001_1100_0011_1000_0001_1100_0011_1000_0001_1100_0011_1000_0001_1100_0011_1000_0001_1100_0011_1111_1111_1100_0011_1111_1111_1100_0011_1111_1111_1100_0011_1000_0001_1100_0011_1000_0001_1100_0011_1000_0001_1100_0011_1000_0001_1100_0011_1000_0001_1100_0000_0000_0000_0000;

localparam S =  256'b0000_0000_0000_0000_0000_1111_1111_1000_0001_1111_1111_1100_0011_1100_0000_0000_0011_1000_0000_0000_0011_1111_0000_0000_0000_1111_1000_0000_0000_1111_1111_0000_0000_0000_1111_1100_0000_0000_0001_1100_0000_0000_0000_1100_0000_0000_0011_1100_0011_1111_1111_0000_0001_1111_1100_0000_0000_0000_0000_0000_0000_0000_0000_0000;

localparam I =  256'b0000_0000_0000_0000_0001_1111_1111_1000_0001_1111_1111_1000_0000_0001_1000_0000_0000_0001_1000_0000_0000_0001_1000_0000_0000_0001_1000_0000_0000_0001_1000_0000_0000_0001_1000_0000_0000_0001_1000_0000_0000_0001_1000_0000_0000_0001_1000_0000_0000_0001_1000_0000_0001_1111_1111_1000_0001_1111_1111_1000_0000_0000_0000_0000;

localparam G =  256'b0000_0000_0000_0000_0000_1111_1111_1000_0000_1111_1111_1100_0011_0000_0000_1100_0011_0000_0000_0000_0011_0000_0000_0000_0011_0000_0000_0000_0011_0000_0000_0000_0011_0000_1111_1000_0011_0000_1111_1100_0011_0000_0000_1100_0011_0000_0000_1100_0011_0000_0000_1100_0000_1111_1111_1100_0000_1111_1111_1000_0000_0000_0000_0000;

localparam N =  256'b0000_0000_0000_0000_0011_1000_0000_1100_0011_1100_0000_1100_0011_1100_0000_1100_0011_1110_0000_1100_0011_0011_0000_1100_0011_0011_0000_1100_0011_0011_0000_1100_0011_0001_1100_1100_0011_0000_1100_1100_0011_0000_1100_1100_0011_0000_0111_1100_0011_0000_0011_1100_0011_0000_0011_1100_0011_0000_0001_1100_0000_0000_0000_0000;

localparam K =  256'b0000_0000_0000_0000_0011_1000_0000_1100_0011_1000_0001_1100_0011_1000_0011_0000_0011_1000_0111_0000_0011_1000_1100_0000_0011_1001_1100_0000_0011_1111_0000_0000_0011_1111_0000_0000_0011_1001_1100_0000_0011_1000_1100_0000_0011_1000_0111_0000_0011_1000_0011_0000_0011_1000_0001_1100_0011_1000_0000_1100_0000_0000_0000_0000;

localparam D =  256'b0000_0000_0000_0000_0011_1111_0000_0000_0011_1111_1100_0000_0011_0000_1111_0000_0011_0000_0111_0000_0011_0000_0001_1000_0011_0000_0001_1000_0011_0000_0000_1100_0011_0000_0000_1100_0011_0000_0001_1000_0011_0000_0001_1000_0011_0000_0111_0000_0011_0000_1111_0000_0011_1111_1100_0000_0011_1111_0000_0000_0000_0000_0000_0000;

localparam P =  256'b0000_0000_0000_0000_0011_1111_1000_0000_0011_1111_1111_0000_0011_0000_0111_1000_0011_0000_0000_1100_0011_0000_0000_1100_0011_0000_0111_1000_0011_1111_1111_0000_0011_1111_1000_0000_0011_0000_0000_0000_0011_0000_0000_0000_0011_0000_0000_0000_0011_0000_0000_0000_0011_0000_0000_0000_0011_0000_0000_0000_0000_0000_0000_0000;

localparam Plus = 256'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001_1000_0000_0000_0001_1000_0000_0000_0001_1000_0000_0000_1111_1111_0000_0000_1111_1111_0000_0000_0001_1000_0000_0000_0001_1000_0000_0000_0001_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;

localparam Minus = 256'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1111_1111_0000_0000_1111_1111_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;

localparam Q =  256'b0000_0000_0000_0000_0000_0011_1100_0000_0000_1111_1111_0000_0001_1100_0011_1000_0011_0000_0000_1100_0011_0000_0000_1100_0011_0000_0000_1100_0011_0000_0000_1100_0011_0000_0000_1100_0011_0000_0000_1100_0011_0000_1100_1100_0011_0000_1110_1100_0001_1100_0111_1000_0000_1111_1111_1100_0000_0011_1100_1100_0000_0000_0000_0000;

localparam T =  256'b0000_0000_0000_0000_0011_1111_1111_1100_0011_1111_1111_1100_0010_0001_1000_0100_0000_0001_1000_0000_0000_0001_1000_0000_0000_0001_1000_0000_0000_0001_1000_0000_0000_0001_1000_0000_0000_0001_1000_0000_0000_0001_1000_0000_0000_0001_1000_0000_0000_0001_1000_0000_0000_0001_1000_0000_0000_0001_1000_0000_0000_0000_0000_0000;

localparam R =  256'b0000_0000_0000_0000_0011_1111_1000_0000_0011_1111_1111_0000_0011_0000_0111_1000_0011_0000_0000_1100_0011_0000_0000_1100_0011_0000_0111_1000_0011_1111_1111_0000_0011_1111_1000_0000_0011_0011_0000_0000_0011_0011_0000_0000_0011_0000_1100_0000_0011_0000_1100_0000_0011_0000_0011_1000_0011_0000_0011_1100_0000_0000_0000_0000;

localparam A =  256'b0000_0000_0000_0000_0000_0111_1110_0000_0000_0111_1110_0000_0000_1100_0011_0000_0001_1100_0011_1000_0011_0000_0000_1100_0011_0000_0000_1100_0011_0000_0000_1100_0011_1111_1111_1100_0011_1111_1111_1100_0011_0000_0000_1100_0011_0000_0000_1100_0011_0000_0000_1100_0011_0000_0000_1100_0011_0000_0000_1100_0000_0000_0000_0000;

//undef
localparam B = 256'b0000_0000_0000_0000_0011_1111_1100_0000_0011_1111_1111_0000_0011_0000_0001_1000_0011_0000_0001_1000_0011_0000_1111_1000_0011_1111_1111_0000_0011_1111_0000_0000_0011_0000_1111_0000_0011_0000_0111_0000_0011_0000_0000_1100_0011_0000_0000_1100_0011_0000_0011_1000_0011_1111_1111_0000_0011_1111_1100_0000_0000_0000_0000_0000;

localparam C = 256'b0000_0000_0000_0000_0000_0111_1111_0000_0001_1111_1111_1000_0011_1000_0000_1100_0011_0000_0000_1100_0011_0000_0000_0000_0011_0000_0000_0000_0011_0000_0000_0000_0011_0000_0000_0000_0011_0000_0000_0000_0011_0000_0000_0000_0011_0000_0000_1100_0011_1000_0000_1100_0001_1111_1111_1000_0000_0111_1111_0000_0000_0000_0000_0000;

localparam E = 256'b0000_0000_0000_0000_0011_1111_1111_1100_0011_1111_1111_1100_0011_0000_0000_1100_0011_0000_0000_1000_0011_0000_0000_0000_0011_0000_0001_0000_0011_1111_1111_0000_0011_1111_1111_0000_0011_0000_0001_0000_0011_0000_0000_0000_0011_0000_0000_1000_0011_0000_0000_1100_0011_1111_1111_1100_0011_1111_1111_1100_0000_0000_0000_0000;

localparam F = 256'b0000_0000_0000_0000_0011_1111_1111_1100_0011_1111_1111_1100_0011_0000_0000_1100_0011_0000_0000_1000_0011_0000_0000_0000_0011_0000_0010_0000_0011_1111_1110_0000_0011_1111_1110_0000_0011_0000_0010_0000_0011_0000_0000_0000_0011_0000_0000_0000_0011_0000_0000_0000_0011_0000_0000_0000_0011_0000_0000_0000_0000_0000_0000_0000;

localparam J = 256'b0000_0000_0000_0000_0011_1111_1111_1100_0011_1111_1111_1100_0000_0001_1000_0000_0000_0001_1000_0000_0000_0001_1000_0000_0000_0001_1000_0000_0000_0001_1000_0000_0000_0001_1000_0000_0000_0001_1000_0000_0000_0001_1000_0000_0010_0001_1000_0000_0011_1001_1000_0000_0011_1111_1000_0000_0000_1111_1000_0000_0000_0000_0000_0000;

localparam L = 256'b0000_0000_0000_0000_0011_0000_0000_0000_0011_0000_0000_0000_0011_0000_0000_0000_0011_0000_0000_0000_0011_0000_0000_0000_0011_0000_0000_0000_0011_0000_0000_0000_0011_0000_0000_0000_0011_0000_0000_0000_0011_0000_0000_0000_0011_0000_0000_0000_0011_0000_0000_0100_0011_1111_1111_1100_0011_1111_1111_1100_0000_0000_0000_0000;

localparam M = 256'b0000_0000_0000_0000_0011_0000_0000_1100_0011_1000_0001_1100_0011_1100_0011_1100_0011_1100_0011_1100_0011_0011_1100_1100_0011_0011_1100_1100_0011_0001_1000_1100_0011_0000_0000_1100_0011_0000_0000_1100_0011_0000_0000_1100_0011_0000_0000_1100_0011_0000_0000_1100_0011_0000_0000_1100_0011_0000_0000_1100_0000_0000_0000_0000;

localparam O = 256'b0000_0000_0000_0000_0000_0011_1100_0000_0000_1111_1111_0000_0001_1100_0011_1000_0011_0000_0000_1100_0011_0000_0000_1100_0011_0000_0000_1100_0011_0000_0000_1100_0011_0000_0000_1100_0011_0000_0000_1100_0011_0000_0000_1100_0011_0000_0000_1100_0001_1100_0011_1000_0000_1111_1111_0000_0000_0011_1100_0000_0000_0000_0000_0000;

localparam U = 256'b0000_0000_0000_0000_0011_0000_0000_1100_0011_0000_0000_1100_0011_0000_0000_1100_0011_0000_0000_1100_0011_0000_0000_1100_0011_0000_0000_1100_0011_0000_0000_1100_0011_0000_0000_1100_0011_0000_0000_1100_0011_0000_0000_1100_0011_0000_0000_1100_0011_0000_0000_1100_0001_1111_1111_1000_0000_1111_1111_0000_0000_0000_0000_0000;

localparam V = 256'b0000_0000_0000_0000_0011_0000_0000_1100_0011_0000_0000_1100_0011_0000_0000_1100_0011_0000_0000_1100_0011_0000_0000_1100_0011_0000_0000_1100_0011_0000_0000_1100_0011_0000_0000_1100_0001_1000_0001_1000_0000_1100_0011_0000_0000_0110_0110_0000_0000_0110_0110_0000_0000_0001_1000_0000_0000_0001_1000_0000_0000_0000_0000_0000;

localparam W = 256'b0000_0000_0000_0000_0011_0000_0000_1100_0011_0000_0000_1100_0011_0000_0000_1100_0011_0000_0000_1100_0011_0000_0000_1100_0011_0000_0000_1100_0011_0000_0000_1100_0011_0000_0000_1100_0011_0001_1000_1100_0011_0001_1000_1100_0011_0011_1100_1100_0011_0011_1100_1100_0001_1100_0011_1000_0000_1100_0011_0000_0000_0000_0000_0000;

localparam X = 256'b0000_0000_0000_0000_0111_0000_0000_1110_0011_0000_0000_1100_0011_0000_0000_1100_0001_1000_0001_1000_0001_1000_0001_1000_0000_1100_0011_0000_0000_1111_1111_0000_0000_1111_1111_0000_0000_1100_0011_0000_0000_1000_0001_0000_0001_1000_0001_1000_0011_0000_0000_1100_0011_0000_0000_1100_0111_0000_0000_1110_0000_0000_0000_0000;

localparam Y = 256'b0000_0000_0000_0000_0111_0000_0000_1110_0011_0000_0000_1100_0011_0000_0000_1100_0001_1000_0001_1000_0001_1100_0011_1000_0000_1110_0111_0000_0000_0111_1110_0000_0000_0001_1000_0000_0000_0001_1000_0000_0000_0001_1000_0000_0000_0001_1000_0000_0000_0001_1000_0000_0000_0001_1000_0000_0000_0001_1000_0000_0000_0000_0000_0000;

localparam Z = 256'b0000_0000_0000_0000_0000_0000_0000_0000_0011_1111_1111_1100_0011_1111_1111_1100_0000_0000_0001_0000_0000_0000_0011_0000_0000_0000_1100_0000_0000_0000_1100_0000_0000_0011_0000_0000_0000_0011_0000_0000_0000_1100_0000_0000_0000_1000_0000_0000_0011_1111_1111_1100_0011_1111_1111_1100_0000_0000_0000_0000_0000_0000_0000_0000;




//

reg [255:0] out;
always @(*) begin 
	case (key)
		8'h16: out = n1; 
		8'h1E: out = n2; 
		8'h26: out = n3; 
		8'h25: out = n4; 
		8'h2E: out = n5; 
		8'h36: out = n6; 
		8'h3D: out = n7; 
		8'h3E: out = n8; 
		8'h46: out = n9; 
		8'h45: out = n0; 
		8'h33: out = H;
		8'h1B: out = S;
		8'h43: out = I;
		8'h34: out = G;
		8'h31: out = N;
		8'h42: out = K;
		8'h23: out = D;
		8'h4D: out = P;
		8'h15: out = Q;
		8'h2C: out = T;
		8'h2D: out = R;
		8'h1C: out = A;
		8'h55: out = Plus;
		8'h4E: out = Minus;
		//undef
		8'h32: out = B;   // b
		8'h21: out = C;   // c
		8'h24: out = E;   // e
		8'h2b: out = F;   // f
		8'h3b: out = J;   // j
		8'h4b: out = L;   // l
		8'h3a: out = M;   // m
		8'h44: out = O;   // o
		8'h3c: out = U;   // u
		8'h2a: out = V;   // v
		8'h1d: out = W;   // w
		8'h22: out = X;   // x
		8'h35: out = Y;   // y
		8'h1a: out = Z;   // z
		8'h0E: out = E;   // show e
		//
		default:
			out = 256'd0;
	endcase 

	o_one_pixel = out[8'd255-{i_Y[4:1], i_X[4:1]}];

end

//1111
//1111
//1111
//1111
//0000
//0000
//0000
//0000
endmodule
